module tb();
  bit a=1'b0;
 
  initial begin
    assert(a)
   
    else
    $warning("The value of a is false");
    
    
  $display("The value of a us %0b",a); 
    
    
  end
 endmodule
